library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity c64rom_basic is
	port (
		clk: in std_logic;
		addr: in unsigned(12 downto 0);
		do: out unsigned(7 downto 0)
	);
end c64rom_basic;

architecture Behavioral of c64rom_basic is
	type romDef is array(0 to  8191) of unsigned(7 downto 0);
	constant romData: romDef := (
		X"94", X"E3", X"7B", X"E3", X"43", X"42", X"4D", X"42", X"41", X"53", X"49", X"43", X"30", X"A8", X"41", X"A7", 
		X"1D", X"AD", X"F7", X"A8", X"A4", X"AB", X"BE", X"AB", X"80", X"B0", X"05", X"AC", X"A4", X"A9", X"9F", X"A8", 
		X"70", X"A8", X"27", X"A9", X"1C", X"A8", X"82", X"A8", X"D1", X"A8", X"3A", X"A9", X"2E", X"A8", X"4A", X"A9", 
		X"2C", X"B8", X"67", X"E1", X"55", X"E1", X"64", X"E1", X"B2", X"B3", X"23", X"B8", X"7F", X"AA", X"9F", X"AA", 
		X"56", X"A8", X"9B", X"A6", X"5D", X"A6", X"85", X"AA", X"29", X"E1", X"BD", X"E1", X"C6", X"E1", X"7A", X"AB", 
		X"41", X"A6", X"39", X"BC", X"CC", X"BC", X"58", X"BC", X"10", X"03", X"7D", X"B3", X"9E", X"B3", X"71", X"BF", 
		X"97", X"E0", X"EA", X"B9", X"ED", X"BF", X"64", X"E2", X"6B", X"E2", X"B4", X"E2", X"0E", X"E3", X"0D", X"B8", 
		X"7C", X"B7", X"65", X"B4", X"AD", X"B7", X"8B", X"B7", X"EC", X"B6", X"00", X"B7", X"2C", X"B7", X"37", X"B7", 
		X"79", X"69", X"B8", X"79", X"52", X"B8", X"7B", X"2A", X"BA", X"7B", X"11", X"BB", X"7F", X"7A", X"BF", X"50", 
		X"E8", X"AF", X"46", X"E5", X"AF", X"7D", X"B3", X"BF", X"5A", X"D3", X"AE", X"64", X"15", X"B0", X"45", X"4E", 
		X"C4", X"46", X"4F", X"D2", X"4E", X"45", X"58", X"D4", X"44", X"41", X"54", X"C1", X"49", X"4E", X"50", X"55", 
		X"54", X"A3", X"49", X"4E", X"50", X"55", X"D4", X"44", X"49", X"CD", X"52", X"45", X"41", X"C4", X"4C", X"45", 
		X"D4", X"47", X"4F", X"54", X"CF", X"52", X"55", X"CE", X"49", X"C6", X"52", X"45", X"53", X"54", X"4F", X"52", 
		X"C5", X"47", X"4F", X"53", X"55", X"C2", X"52", X"45", X"54", X"55", X"52", X"CE", X"52", X"45", X"CD", X"53", 
		X"54", X"4F", X"D0", X"4F", X"CE", X"57", X"41", X"49", X"D4", X"4C", X"4F", X"41", X"C4", X"53", X"41", X"56", 
		X"C5", X"56", X"45", X"52", X"49", X"46", X"D9", X"44", X"45", X"C6", X"50", X"4F", X"4B", X"C5", X"50", X"52", 
		X"49", X"4E", X"54", X"A3", X"50", X"52", X"49", X"4E", X"D4", X"43", X"4F", X"4E", X"D4", X"4C", X"49", X"53", 
		X"D4", X"43", X"4C", X"D2", X"43", X"4D", X"C4", X"53", X"59", X"D3", X"4F", X"50", X"45", X"CE", X"43", X"4C", 
		X"4F", X"53", X"C5", X"47", X"45", X"D4", X"4E", X"45", X"D7", X"54", X"41", X"42", X"A8", X"54", X"CF", X"46", 
		X"CE", X"53", X"50", X"43", X"A8", X"54", X"48", X"45", X"CE", X"4E", X"4F", X"D4", X"53", X"54", X"45", X"D0", 
		X"AB", X"AD", X"AA", X"AF", X"DE", X"41", X"4E", X"C4", X"4F", X"D2", X"BE", X"BD", X"BC", X"53", X"47", X"CE", 
		X"49", X"4E", X"D4", X"41", X"42", X"D3", X"55", X"53", X"D2", X"46", X"52", X"C5", X"50", X"4F", X"D3", X"53", 
		X"51", X"D2", X"52", X"4E", X"C4", X"4C", X"4F", X"C7", X"45", X"58", X"D0", X"43", X"4F", X"D3", X"53", X"49", 
		X"CE", X"54", X"41", X"CE", X"41", X"54", X"CE", X"50", X"45", X"45", X"CB", X"4C", X"45", X"CE", X"53", X"54", 
		X"52", X"A4", X"56", X"41", X"CC", X"41", X"53", X"C3", X"43", X"48", X"52", X"A4", X"4C", X"45", X"46", X"54", 
		X"A4", X"52", X"49", X"47", X"48", X"54", X"A4", X"4D", X"49", X"44", X"A4", X"47", X"CF", X"00", X"54", X"4F", 
		X"4F", X"20", X"4D", X"41", X"4E", X"59", X"20", X"46", X"49", X"4C", X"45", X"D3", X"46", X"49", X"4C", X"45", 
		X"20", X"4F", X"50", X"45", X"CE", X"46", X"49", X"4C", X"45", X"20", X"4E", X"4F", X"54", X"20", X"4F", X"50", 
		X"45", X"CE", X"46", X"49", X"4C", X"45", X"20", X"4E", X"4F", X"54", X"20", X"46", X"4F", X"55", X"4E", X"C4", 
		X"44", X"45", X"56", X"49", X"43", X"45", X"20", X"4E", X"4F", X"54", X"20", X"50", X"52", X"45", X"53", X"45", 
		X"4E", X"D4", X"4E", X"4F", X"54", X"20", X"49", X"4E", X"50", X"55", X"54", X"20", X"46", X"49", X"4C", X"C5", 
		X"4E", X"4F", X"54", X"20", X"4F", X"55", X"54", X"50", X"55", X"54", X"20", X"46", X"49", X"4C", X"C5", X"4D", 
		X"49", X"53", X"53", X"49", X"4E", X"47", X"20", X"46", X"49", X"4C", X"45", X"20", X"4E", X"41", X"4D", X"C5", 
		X"49", X"4C", X"4C", X"45", X"47", X"41", X"4C", X"20", X"44", X"45", X"56", X"49", X"43", X"45", X"20", X"4E", 
		X"55", X"4D", X"42", X"45", X"D2", X"4E", X"45", X"58", X"54", X"20", X"57", X"49", X"54", X"48", X"4F", X"55", 
		X"54", X"20", X"46", X"4F", X"D2", X"53", X"59", X"4E", X"54", X"41", X"D8", X"52", X"45", X"54", X"55", X"52", 
		X"4E", X"20", X"57", X"49", X"54", X"48", X"4F", X"55", X"54", X"20", X"47", X"4F", X"53", X"55", X"C2", X"4F", 
		X"55", X"54", X"20", X"4F", X"46", X"20", X"44", X"41", X"54", X"C1", X"49", X"4C", X"4C", X"45", X"47", X"41", 
		X"4C", X"20", X"51", X"55", X"41", X"4E", X"54", X"49", X"54", X"D9", X"4F", X"56", X"45", X"52", X"46", X"4C", 
		X"4F", X"D7", X"4F", X"55", X"54", X"20", X"4F", X"46", X"20", X"4D", X"45", X"4D", X"4F", X"52", X"D9", X"55", 
		X"4E", X"44", X"45", X"46", X"27", X"44", X"20", X"53", X"54", X"41", X"54", X"45", X"4D", X"45", X"4E", X"D4", 
		X"42", X"41", X"44", X"20", X"53", X"55", X"42", X"53", X"43", X"52", X"49", X"50", X"D4", X"52", X"45", X"44", 
		X"49", X"4D", X"27", X"44", X"20", X"41", X"52", X"52", X"41", X"D9", X"44", X"49", X"56", X"49", X"53", X"49", 
		X"4F", X"4E", X"20", X"42", X"59", X"20", X"5A", X"45", X"52", X"CF", X"49", X"4C", X"4C", X"45", X"47", X"41", 
		X"4C", X"20", X"44", X"49", X"52", X"45", X"43", X"D4", X"54", X"59", X"50", X"45", X"20", X"4D", X"49", X"53", 
		X"4D", X"41", X"54", X"43", X"C8", X"53", X"54", X"52", X"49", X"4E", X"47", X"20", X"54", X"4F", X"4F", X"20", 
		X"4C", X"4F", X"4E", X"C7", X"46", X"49", X"4C", X"45", X"20", X"44", X"41", X"54", X"C1", X"46", X"4F", X"52", 
		X"4D", X"55", X"4C", X"41", X"20", X"54", X"4F", X"4F", X"20", X"43", X"4F", X"4D", X"50", X"4C", X"45", X"D8", 
		X"43", X"41", X"4E", X"27", X"54", X"20", X"43", X"4F", X"4E", X"54", X"49", X"4E", X"55", X"C5", X"55", X"4E", 
		X"44", X"45", X"46", X"27", X"44", X"20", X"46", X"55", X"4E", X"43", X"54", X"49", X"4F", X"CE", X"56", X"45", 
		X"52", X"49", X"46", X"D9", X"4C", X"4F", X"41", X"C4", X"9E", X"A1", X"AC", X"A1", X"B5", X"A1", X"C2", X"A1", 
		X"D0", X"A1", X"E2", X"A1", X"F0", X"A1", X"FF", X"A1", X"10", X"A2", X"25", X"A2", X"35", X"A2", X"3B", X"A2", 
		X"4F", X"A2", X"5A", X"A2", X"6A", X"A2", X"72", X"A2", X"7F", X"A2", X"90", X"A2", X"9D", X"A2", X"AA", X"A2", 
		X"BA", X"A2", X"C8", X"A2", X"D5", X"A2", X"E4", X"A2", X"ED", X"A2", X"00", X"A3", X"0E", X"A3", X"1E", X"A3", 
		X"24", X"A3", X"83", X"A3", X"0D", X"4F", X"4B", X"0D", X"00", X"20", X"20", X"45", X"52", X"52", X"4F", X"52", 
		X"00", X"20", X"49", X"4E", X"20", X"00", X"0D", X"0A", X"52", X"45", X"41", X"44", X"59", X"2E", X"0D", X"0A", 
		X"00", X"0D", X"0A", X"42", X"52", X"45", X"41", X"4B", X"00", X"A0", X"BA", X"E8", X"E8", X"E8", X"E8", X"BD", 
		X"01", X"01", X"C9", X"81", X"D0", X"21", X"A5", X"4A", X"D0", X"0A", X"BD", X"02", X"01", X"85", X"49", X"BD", 
		X"03", X"01", X"85", X"4A", X"DD", X"03", X"01", X"D0", X"07", X"A5", X"49", X"DD", X"02", X"01", X"F0", X"07", 
		X"8A", X"18", X"69", X"12", X"AA", X"D0", X"D8", X"60", X"20", X"08", X"A4", X"85", X"31", X"84", X"32", X"38", 
		X"A5", X"5A", X"E5", X"5F", X"85", X"22", X"A8", X"A5", X"5B", X"E5", X"60", X"AA", X"E8", X"98", X"F0", X"23", 
		X"A5", X"5A", X"38", X"E5", X"22", X"85", X"5A", X"B0", X"03", X"C6", X"5B", X"38", X"A5", X"58", X"E5", X"22", 
		X"85", X"58", X"B0", X"08", X"C6", X"59", X"90", X"04", X"B1", X"5A", X"91", X"58", X"88", X"D0", X"F9", X"B1", 
		X"5A", X"91", X"58", X"C6", X"5B", X"C6", X"59", X"CA", X"D0", X"F2", X"60", X"0A", X"69", X"3E", X"B0", X"35", 
		X"85", X"22", X"BA", X"E4", X"22", X"90", X"2E", X"60", X"C4", X"34", X"90", X"28", X"D0", X"04", X"C5", X"33", 
		X"90", X"22", X"48", X"A2", X"09", X"98", X"48", X"B5", X"57", X"CA", X"10", X"FA", X"20", X"26", X"B5", X"A2", 
		X"F7", X"68", X"95", X"61", X"E8", X"30", X"FA", X"68", X"A8", X"68", X"C4", X"34", X"90", X"06", X"D0", X"05", 
		X"C5", X"33", X"B0", X"01", X"60", X"A2", X"10", X"6C", X"00", X"03", X"8A", X"0A", X"AA", X"BD", X"26", X"A3", 
		X"85", X"22", X"BD", X"27", X"A3", X"85", X"23", X"20", X"CC", X"FF", X"A9", X"00", X"85", X"13", X"20", X"D7", 
		X"AA", X"20", X"45", X"AB", X"A0", X"00", X"B1", X"22", X"48", X"29", X"7F", X"20", X"47", X"AB", X"C8", X"68", 
		X"10", X"F4", X"20", X"7A", X"A6", X"A9", X"69", X"A0", X"A3", X"20", X"1E", X"AB", X"A4", X"3A", X"C8", X"F0", 
		X"03", X"20", X"C2", X"BD", X"A9", X"76", X"A0", X"A3", X"20", X"1E", X"AB", X"A9", X"80", X"20", X"90", X"FF", 
		X"6C", X"02", X"03", X"20", X"60", X"A5", X"86", X"7A", X"84", X"7B", X"20", X"73", X"00", X"AA", X"F0", X"F0", 
		X"A2", X"FF", X"86", X"3A", X"90", X"06", X"20", X"79", X"A5", X"4C", X"E1", X"A7", X"20", X"6B", X"A9", X"20", 
		X"79", X"A5", X"84", X"0B", X"20", X"13", X"A6", X"90", X"44", X"A0", X"01", X"B1", X"5F", X"85", X"23", X"A5", 
		X"2D", X"85", X"22", X"A5", X"60", X"85", X"25", X"A5", X"5F", X"88", X"F1", X"5F", X"18", X"65", X"2D", X"85", 
		X"2D", X"85", X"24", X"A5", X"2E", X"69", X"FF", X"85", X"2E", X"E5", X"60", X"AA", X"38", X"A5", X"5F", X"E5", 
		X"2D", X"A8", X"B0", X"03", X"E8", X"C6", X"25", X"18", X"65", X"22", X"90", X"03", X"C6", X"23", X"18", X"B1", 
		X"22", X"91", X"24", X"C8", X"D0", X"F9", X"E6", X"23", X"E6", X"25", X"CA", X"D0", X"F2", X"20", X"59", X"A6", 
		X"20", X"33", X"A5", X"AD", X"00", X"02", X"F0", X"88", X"18", X"A5", X"2D", X"85", X"5A", X"65", X"0B", X"85", 
		X"58", X"A4", X"2E", X"84", X"5B", X"90", X"01", X"C8", X"84", X"59", X"20", X"B8", X"A3", X"A5", X"14", X"A4", 
		X"15", X"8D", X"FE", X"01", X"8C", X"FF", X"01", X"A5", X"31", X"A4", X"32", X"85", X"2D", X"84", X"2E", X"A4", 
		X"0B", X"88", X"B9", X"FC", X"01", X"91", X"5F", X"88", X"10", X"F8", X"20", X"59", X"A6", X"20", X"33", X"A5", 
		X"4C", X"80", X"A4", X"A5", X"2B", X"A4", X"2C", X"85", X"22", X"84", X"23", X"18", X"A0", X"01", X"B1", X"22", 
		X"F0", X"1D", X"A0", X"04", X"C8", X"B1", X"22", X"D0", X"FB", X"C8", X"98", X"65", X"22", X"AA", X"A0", X"00", 
		X"91", X"22", X"A5", X"23", X"69", X"00", X"C8", X"91", X"22", X"86", X"22", X"85", X"23", X"90", X"DD", X"60", 
		X"A2", X"00", X"20", X"12", X"E1", X"C9", X"0D", X"F0", X"0D", X"9D", X"00", X"02", X"E8", X"E0", X"59", X"90", 
		X"F1", X"A2", X"17", X"4C", X"37", X"A4", X"4C", X"CA", X"AA", X"6C", X"04", X"03", X"A6", X"7A", X"A0", X"04", 
		X"84", X"0F", X"BD", X"00", X"02", X"10", X"07", X"C9", X"FF", X"F0", X"3E", X"E8", X"D0", X"F4", X"C9", X"20", 
		X"F0", X"37", X"85", X"08", X"C9", X"22", X"F0", X"56", X"24", X"0F", X"70", X"2D", X"C9", X"3F", X"D0", X"04", 
		X"A9", X"99", X"D0", X"25", X"C9", X"30", X"90", X"04", X"C9", X"3C", X"90", X"1D", X"84", X"71", X"A0", X"00", 
		X"84", X"0B", X"88", X"86", X"7A", X"CA", X"C8", X"E8", X"BD", X"00", X"02", X"38", X"F9", X"9E", X"A0", X"F0", 
		X"F5", X"C9", X"80", X"D0", X"30", X"05", X"0B", X"A4", X"71", X"E8", X"C8", X"99", X"FB", X"01", X"B9", X"FB", 
		X"01", X"F0", X"36", X"38", X"E9", X"3A", X"F0", X"04", X"C9", X"49", X"D0", X"02", X"85", X"0F", X"38", X"E9", 
		X"55", X"D0", X"9F", X"85", X"08", X"BD", X"00", X"02", X"F0", X"DF", X"C5", X"08", X"F0", X"DB", X"C8", X"99", 
		X"FB", X"01", X"E8", X"D0", X"F0", X"A6", X"7A", X"E6", X"0B", X"C8", X"B9", X"9D", X"A0", X"10", X"FA", X"B9", 
		X"9E", X"A0", X"D0", X"B4", X"BD", X"00", X"02", X"10", X"BE", X"99", X"FD", X"01", X"C6", X"7B", X"A9", X"FF", 
		X"85", X"7A", X"60", X"A5", X"2B", X"A6", X"2C", X"A0", X"01", X"85", X"5F", X"86", X"60", X"B1", X"5F", X"F0", 
		X"1F", X"C8", X"C8", X"A5", X"15", X"D1", X"5F", X"90", X"18", X"F0", X"03", X"88", X"D0", X"09", X"A5", X"14", 
		X"88", X"D1", X"5F", X"90", X"0C", X"F0", X"0A", X"88", X"B1", X"5F", X"AA", X"88", X"B1", X"5F", X"B0", X"D7", 
		X"18", X"60", X"D0", X"FD", X"A9", X"00", X"A8", X"91", X"2B", X"C8", X"91", X"2B", X"A5", X"2B", X"18", X"69", 
		X"02", X"85", X"2D", X"A5", X"2C", X"69", X"00", X"85", X"2E", X"20", X"8E", X"A6", X"A9", X"00", X"D0", X"2D", 
		X"20", X"E7", X"FF", X"A5", X"37", X"A4", X"38", X"85", X"33", X"84", X"34", X"A5", X"2D", X"A4", X"2E", X"85", 
		X"2F", X"84", X"30", X"85", X"31", X"84", X"32", X"20", X"1D", X"A8", X"A2", X"19", X"86", X"16", X"68", X"A8", 
		X"68", X"A2", X"FA", X"9A", X"48", X"98", X"48", X"A9", X"00", X"85", X"3E", X"85", X"10", X"60", X"18", X"A5", 
		X"2B", X"69", X"FF", X"85", X"7A", X"A5", X"2C", X"69", X"FF", X"85", X"7B", X"60", X"90", X"06", X"F0", X"04", 
		X"C9", X"AB", X"D0", X"E9", X"20", X"6B", X"A9", X"20", X"13", X"A6", X"20", X"79", X"00", X"F0", X"0C", X"C9", 
		X"AB", X"D0", X"8E", X"20", X"73", X"00", X"20", X"6B", X"A9", X"D0", X"86", X"68", X"68", X"A5", X"14", X"05", 
		X"15", X"D0", X"06", X"A9", X"FF", X"85", X"14", X"85", X"15", X"A0", X"01", X"84", X"0F", X"B1", X"5F", X"F0", 
		X"43", X"20", X"2C", X"A8", X"20", X"D7", X"AA", X"C8", X"B1", X"5F", X"AA", X"C8", X"B1", X"5F", X"C5", X"15", 
		X"D0", X"04", X"E4", X"14", X"F0", X"02", X"B0", X"2C", X"84", X"49", X"20", X"CD", X"BD", X"A9", X"20", X"A4", 
		X"49", X"29", X"7F", X"20", X"47", X"AB", X"C9", X"22", X"D0", X"06", X"A5", X"0F", X"49", X"FF", X"85", X"0F", 
		X"C8", X"F0", X"11", X"B1", X"5F", X"D0", X"10", X"A8", X"B1", X"5F", X"AA", X"C8", X"B1", X"5F", X"86", X"5F", 
		X"85", X"60", X"D0", X"B5", X"4C", X"86", X"E3", X"6C", X"06", X"03", X"10", X"D7", X"C9", X"FF", X"F0", X"D3", 
		X"24", X"0F", X"30", X"CF", X"38", X"E9", X"7F", X"AA", X"84", X"49", X"A0", X"FF", X"CA", X"F0", X"08", X"C8", 
		X"B9", X"9E", X"A0", X"10", X"FA", X"30", X"F5", X"C8", X"B9", X"9E", X"A0", X"30", X"B2", X"20", X"47", X"AB", 
		X"D0", X"F5", X"A9", X"80", X"85", X"10", X"20", X"A5", X"A9", X"20", X"8A", X"A3", X"D0", X"05", X"8A", X"69", 
		X"0F", X"AA", X"9A", X"68", X"68", X"A9", X"09", X"20", X"FB", X"A3", X"20", X"06", X"A9", X"18", X"98", X"65", 
		X"7A", X"48", X"A5", X"7B", X"69", X"00", X"48", X"A5", X"3A", X"48", X"A5", X"39", X"48", X"A9", X"A4", X"20", 
		X"FF", X"AE", X"20", X"8D", X"AD", X"20", X"8A", X"AD", X"A5", X"66", X"09", X"7F", X"25", X"62", X"85", X"62", 
		X"A9", X"8B", X"A0", X"A7", X"85", X"22", X"84", X"23", X"4C", X"43", X"AE", X"A9", X"BC", X"A0", X"B9", X"20", 
		X"A2", X"BB", X"20", X"79", X"00", X"C9", X"A9", X"D0", X"06", X"20", X"73", X"00", X"20", X"8A", X"AD", X"20", 
		X"2B", X"BC", X"20", X"38", X"AE", X"A5", X"4A", X"48", X"A5", X"49", X"48", X"A9", X"81", X"48", X"20", X"2C", 
		X"A8", X"A5", X"7A", X"A4", X"7B", X"C0", X"02", X"EA", X"F0", X"04", X"85", X"3D", X"84", X"3E", X"A0", X"00", 
		X"B1", X"7A", X"D0", X"43", X"A0", X"02", X"B1", X"7A", X"18", X"D0", X"03", X"4C", X"4B", X"A8", X"C8", X"B1", 
		X"7A", X"85", X"39", X"C8", X"B1", X"7A", X"85", X"3A", X"98", X"65", X"7A", X"85", X"7A", X"90", X"02", X"E6", 
		X"7B", X"6C", X"08", X"03", X"20", X"73", X"00", X"20", X"ED", X"A7", X"4C", X"AE", X"A7", X"F0", X"3C", X"E9", 
		X"80", X"90", X"11", X"C9", X"23", X"B0", X"17", X"0A", X"A8", X"B9", X"0D", X"A0", X"48", X"B9", X"0C", X"A0", 
		X"48", X"4C", X"73", X"00", X"4C", X"A5", X"A9", X"C9", X"3A", X"F0", X"D6", X"4C", X"08", X"AF", X"C9", X"4B", 
		X"D0", X"F9", X"20", X"73", X"00", X"A9", X"A4", X"20", X"FF", X"AE", X"4C", X"A0", X"A8", X"38", X"A5", X"2B", 
		X"E9", X"01", X"A4", X"2C", X"B0", X"01", X"88", X"85", X"41", X"84", X"42", X"60", X"20", X"E1", X"FF", X"B0", 
		X"01", X"18", X"D0", X"3C", X"A5", X"7A", X"A4", X"7B", X"A6", X"3A", X"E8", X"F0", X"0C", X"85", X"3D", X"84", 
		X"3E", X"A5", X"39", X"A4", X"3A", X"85", X"3B", X"84", X"3C", X"68", X"68", X"A9", X"81", X"A0", X"A3", X"90", 
		X"03", X"4C", X"69", X"A4", X"4C", X"86", X"E3", X"D0", X"17", X"A2", X"1A", X"A4", X"3E", X"D0", X"03", X"4C", 
		X"37", X"A4", X"A5", X"3D", X"85", X"7A", X"84", X"7B", X"A5", X"3B", X"A4", X"3C", X"85", X"39", X"84", X"3A", 
		X"60", X"08", X"A9", X"00", X"20", X"90", X"FF", X"28", X"D0", X"03", X"4C", X"59", X"A6", X"20", X"60", X"A6", 
		X"4C", X"97", X"A8", X"A9", X"03", X"20", X"FB", X"A3", X"A5", X"7B", X"48", X"A5", X"7A", X"48", X"A5", X"3A", 
		X"48", X"A5", X"39", X"48", X"A9", X"8D", X"48", X"20", X"79", X"00", X"20", X"A0", X"A8", X"4C", X"AE", X"A7", 
		X"20", X"6B", X"A9", X"20", X"09", X"A9", X"38", X"A5", X"39", X"E5", X"14", X"A5", X"3A", X"E5", X"15", X"B0", 
		X"0B", X"98", X"38", X"65", X"7A", X"A6", X"7B", X"90", X"07", X"E8", X"B0", X"04", X"A5", X"2B", X"A6", X"2C", 
		X"20", X"17", X"A6", X"90", X"1E", X"A5", X"5F", X"E9", X"01", X"85", X"7A", X"A5", X"60", X"E9", X"00", X"85", 
		X"7B", X"60", X"D0", X"FD", X"A9", X"FF", X"85", X"4A", X"20", X"8A", X"A3", X"9A", X"C9", X"8D", X"F0", X"0B", 
		X"A2", X"0C", X"2C", X"A2", X"11", X"4C", X"37", X"A4", X"4C", X"08", X"AF", X"68", X"68", X"85", X"39", X"68", 
		X"85", X"3A", X"68", X"85", X"7A", X"68", X"85", X"7B", X"20", X"06", X"A9", X"98", X"18", X"65", X"7A", X"85", 
		X"7A", X"90", X"02", X"E6", X"7B", X"60", X"A2", X"3A", X"2C", X"A2", X"00", X"86", X"07", X"A0", X"00", X"84", 
		X"08", X"A5", X"08", X"A6", X"07", X"85", X"07", X"86", X"08", X"B1", X"7A", X"F0", X"E8", X"C5", X"08", X"F0", 
		X"E4", X"C8", X"C9", X"22", X"D0", X"F3", X"F0", X"E9", X"20", X"9E", X"AD", X"20", X"79", X"00", X"C9", X"89", 
		X"F0", X"05", X"A9", X"A7", X"20", X"FF", X"AE", X"A5", X"61", X"D0", X"05", X"20", X"09", X"A9", X"F0", X"BB", 
		X"20", X"79", X"00", X"B0", X"03", X"4C", X"A0", X"A8", X"4C", X"ED", X"A7", X"20", X"9E", X"B7", X"48", X"C9", 
		X"8D", X"F0", X"04", X"C9", X"89", X"D0", X"91", X"C6", X"65", X"D0", X"04", X"68", X"4C", X"EF", X"A7", X"20", 
		X"73", X"00", X"20", X"6B", X"A9", X"C9", X"2C", X"F0", X"EE", X"68", X"60", X"A2", X"00", X"86", X"14", X"86", 
		X"15", X"B0", X"F7", X"E9", X"2F", X"85", X"07", X"A5", X"15", X"85", X"22", X"C9", X"19", X"B0", X"D4", X"A5", 
		X"14", X"0A", X"26", X"22", X"0A", X"26", X"22", X"65", X"14", X"85", X"14", X"A5", X"22", X"65", X"15", X"85", 
		X"15", X"06", X"14", X"26", X"15", X"A5", X"14", X"65", X"07", X"85", X"14", X"90", X"02", X"E6", X"15", X"20", 
		X"73", X"00", X"4C", X"71", X"A9", X"20", X"8B", X"B0", X"85", X"49", X"84", X"4A", X"A9", X"B2", X"20", X"FF", 
		X"AE", X"A5", X"0E", X"48", X"A5", X"0D", X"48", X"20", X"9E", X"AD", X"68", X"2A", X"20", X"90", X"AD", X"D0", 
		X"18", X"68", X"10", X"12", X"20", X"1B", X"BC", X"20", X"BF", X"B1", X"A0", X"00", X"A5", X"64", X"91", X"49", 
		X"C8", X"A5", X"65", X"91", X"49", X"60", X"4C", X"D0", X"BB", X"68", X"A4", X"4A", X"C0", X"BF", X"D0", X"4C", 
		X"20", X"A6", X"B6", X"C9", X"06", X"D0", X"3D", X"A0", X"00", X"84", X"61", X"84", X"66", X"84", X"71", X"20", 
		X"1D", X"AA", X"20", X"E2", X"BA", X"E6", X"71", X"A4", X"71", X"20", X"1D", X"AA", X"20", X"0C", X"BC", X"AA", 
		X"F0", X"05", X"E8", X"8A", X"20", X"ED", X"BA", X"A4", X"71", X"C8", X"C0", X"06", X"D0", X"DF", X"20", X"E2", 
		X"BA", X"20", X"9B", X"BC", X"A6", X"64", X"A4", X"63", X"A5", X"65", X"4C", X"DB", X"FF", X"B1", X"22", X"20", 
		X"80", X"00", X"90", X"03", X"4C", X"48", X"B2", X"E9", X"2F", X"4C", X"7E", X"BD", X"A0", X"02", X"B1", X"64", 
		X"C5", X"34", X"90", X"17", X"D0", X"07", X"88", X"B1", X"64", X"C5", X"33", X"90", X"0E", X"A4", X"65", X"C4", 
		X"2E", X"90", X"08", X"D0", X"0D", X"A5", X"64", X"C5", X"2D", X"B0", X"07", X"A5", X"64", X"A4", X"65", X"4C", 
		X"68", X"AA", X"A0", X"00", X"B1", X"64", X"20", X"75", X"B4", X"A5", X"50", X"A4", X"51", X"85", X"6F", X"84", 
		X"70", X"20", X"7A", X"B6", X"A9", X"61", X"A0", X"00", X"85", X"50", X"84", X"51", X"20", X"DB", X"B6", X"A0", 
		X"00", X"B1", X"50", X"91", X"49", X"C8", X"B1", X"50", X"91", X"49", X"C8", X"B1", X"50", X"91", X"49", X"60", 
		X"20", X"86", X"AA", X"4C", X"B5", X"AB", X"20", X"9E", X"B7", X"F0", X"05", X"A9", X"2C", X"20", X"FF", X"AE", 
		X"08", X"86", X"13", X"20", X"18", X"E1", X"28", X"4C", X"A0", X"AA", X"20", X"21", X"AB", X"20", X"79", X"00", 
		X"F0", X"35", X"F0", X"43", X"C9", X"A3", X"F0", X"50", X"C9", X"A6", X"18", X"F0", X"4B", X"C9", X"2C", X"F0", 
		X"37", X"C9", X"3B", X"F0", X"5E", X"20", X"9E", X"AD", X"24", X"0D", X"30", X"DE", X"20", X"DD", X"BD", X"20", 
		X"87", X"B4", X"20", X"21", X"AB", X"20", X"3B", X"AB", X"D0", X"D3", X"A9", X"00", X"9D", X"00", X"02", X"A2", 
		X"FF", X"A0", X"01", X"A5", X"13", X"D0", X"10", X"A9", X"0D", X"20", X"47", X"AB", X"24", X"13", X"10", X"05", 
		X"A9", X"0A", X"20", X"47", X"AB", X"49", X"FF", X"60", X"38", X"20", X"F0", X"FF", X"98", X"38", X"E9", X"0A", 
		X"B0", X"FC", X"49", X"FF", X"69", X"01", X"D0", X"16", X"08", X"38", X"20", X"F0", X"FF", X"84", X"09", X"20", 
		X"9B", X"B7", X"C9", X"29", X"D0", X"59", X"28", X"90", X"06", X"8A", X"E5", X"09", X"90", X"05", X"AA", X"E8", 
		X"CA", X"D0", X"06", X"20", X"73", X"00", X"4C", X"A2", X"AA", X"20", X"3B", X"AB", X"D0", X"F2", X"20", X"87", 
		X"B4", X"20", X"A6", X"B6", X"AA", X"A0", X"00", X"E8", X"CA", X"F0", X"BC", X"B1", X"22", X"20", X"47", X"AB", 
		X"C8", X"C9", X"0D", X"D0", X"F3", X"20", X"E5", X"AA", X"4C", X"28", X"AB", X"A5", X"13", X"F0", X"03", X"A9", 
		X"20", X"2C", X"A9", X"1D", X"2C", X"A9", X"3F", X"20", X"0C", X"E1", X"29", X"FF", X"60", X"A5", X"11", X"F0", 
		X"11", X"30", X"04", X"A0", X"FF", X"D0", X"04", X"A5", X"3F", X"A4", X"40", X"85", X"39", X"84", X"3A", X"4C", 
		X"08", X"AF", X"A5", X"13", X"F0", X"05", X"A2", X"18", X"4C", X"37", X"A4", X"A9", X"0C", X"A0", X"AD", X"20", 
		X"1E", X"AB", X"A5", X"3D", X"A4", X"3E", X"85", X"7A", X"84", X"7B", X"60", X"20", X"A6", X"B3", X"C9", X"23", 
		X"D0", X"10", X"20", X"73", X"00", X"20", X"9E", X"B7", X"A9", X"2C", X"20", X"FF", X"AE", X"86", X"13", X"20", 
		X"1E", X"E1", X"A2", X"01", X"A0", X"02", X"A9", X"00", X"8D", X"01", X"02", X"A9", X"40", X"20", X"0F", X"AC", 
		X"A6", X"13", X"D0", X"13", X"60", X"20", X"9E", X"B7", X"A9", X"2C", X"20", X"FF", X"AE", X"86", X"13", X"20", 
		X"1E", X"E1", X"20", X"CE", X"AB", X"A5", X"13", X"20", X"CC", X"FF", X"A2", X"00", X"86", X"13", X"60", X"C9", 
		X"22", X"D0", X"0B", X"20", X"BD", X"AE", X"A9", X"3B", X"20", X"FF", X"AE", X"20", X"21", X"AB", X"20", X"A6", 
		X"B3", X"A9", X"2C", X"8D", X"FF", X"01", X"20", X"F9", X"AB", X"A5", X"13", X"F0", X"0D", X"20", X"B7", X"FF", 
		X"29", X"02", X"F0", X"06", X"20", X"B5", X"AB", X"4C", X"F8", X"A8", X"AD", X"00", X"02", X"D0", X"1E", X"A5", 
		X"13", X"D0", X"E3", X"20", X"06", X"A9", X"4C", X"FB", X"A8", X"A5", X"13", X"D0", X"06", X"20", X"45", X"AB", 
		X"20", X"3B", X"AB", X"4C", X"60", X"A5", X"A6", X"41", X"A4", X"42", X"A9", X"98", X"2C", X"A9", X"00", X"85", 
		X"11", X"86", X"43", X"84", X"44", X"20", X"8B", X"B0", X"85", X"49", X"84", X"4A", X"A5", X"7A", X"A4", X"7B", 
		X"85", X"4B", X"84", X"4C", X"A6", X"43", X"A4", X"44", X"86", X"7A", X"84", X"7B", X"20", X"79", X"00", X"D0", 
		X"20", X"24", X"11", X"50", X"0C", X"20", X"24", X"E1", X"8D", X"00", X"02", X"A2", X"FF", X"A0", X"01", X"D0", 
		X"0C", X"30", X"75", X"A5", X"13", X"D0", X"03", X"20", X"45", X"AB", X"20", X"F9", X"AB", X"86", X"7A", X"84", 
		X"7B", X"20", X"73", X"00", X"24", X"0D", X"10", X"31", X"24", X"11", X"50", X"09", X"E8", X"86", X"7A", X"A9", 
		X"00", X"85", X"07", X"F0", X"0C", X"85", X"07", X"C9", X"22", X"F0", X"07", X"A9", X"3A", X"85", X"07", X"A9", 
		X"2C", X"18", X"85", X"08", X"A5", X"7A", X"A4", X"7B", X"69", X"00", X"90", X"01", X"C8", X"20", X"8D", X"B4", 
		X"20", X"E2", X"B7", X"20", X"DA", X"A9", X"4C", X"91", X"AC", X"20", X"F3", X"BC", X"A5", X"0E", X"20", X"C2", 
		X"A9", X"20", X"79", X"00", X"F0", X"07", X"C9", X"2C", X"F0", X"03", X"4C", X"4D", X"AB", X"A5", X"7A", X"A4", 
		X"7B", X"85", X"43", X"84", X"44", X"A5", X"4B", X"A4", X"4C", X"85", X"7A", X"84", X"7B", X"20", X"79", X"00", 
		X"F0", X"2D", X"20", X"FD", X"AE", X"4C", X"15", X"AC", X"20", X"06", X"A9", X"C8", X"AA", X"D0", X"12", X"A2", 
		X"0D", X"C8", X"B1", X"7A", X"F0", X"6C", X"C8", X"B1", X"7A", X"85", X"3F", X"C8", X"B1", X"7A", X"C8", X"85", 
		X"40", X"20", X"FB", X"A8", X"20", X"79", X"00", X"AA", X"E0", X"83", X"D0", X"DC", X"4C", X"51", X"AC", X"A5", 
		X"43", X"A4", X"44", X"A6", X"11", X"10", X"03", X"4C", X"27", X"A8", X"A0", X"00", X"B1", X"43", X"F0", X"0B", 
		X"A5", X"13", X"D0", X"07", X"A9", X"FC", X"A0", X"AC", X"4C", X"1E", X"AB", X"60", X"3F", X"45", X"58", X"54", 
		X"52", X"41", X"20", X"49", X"47", X"4E", X"4F", X"52", X"45", X"44", X"0D", X"00", X"3F", X"52", X"45", X"44", 
		X"4F", X"20", X"46", X"52", X"4F", X"4D", X"20", X"53", X"54", X"41", X"52", X"54", X"0D", X"00", X"D0", X"04", 
		X"A0", X"00", X"F0", X"03", X"20", X"8B", X"B0", X"85", X"49", X"84", X"4A", X"20", X"8A", X"A3", X"F0", X"05", 
		X"A2", X"0A", X"4C", X"37", X"A4", X"9A", X"8A", X"18", X"69", X"04", X"48", X"69", X"06", X"85", X"24", X"68", 
		X"A0", X"01", X"20", X"A2", X"BB", X"BA", X"BD", X"09", X"01", X"85", X"66", X"A5", X"49", X"A4", X"4A", X"20", 
		X"67", X"B8", X"20", X"D0", X"BB", X"A0", X"01", X"20", X"5D", X"BC", X"BA", X"38", X"FD", X"09", X"01", X"F0", 
		X"17", X"BD", X"0F", X"01", X"85", X"39", X"BD", X"10", X"01", X"85", X"3A", X"BD", X"12", X"01", X"85", X"7A", 
		X"BD", X"11", X"01", X"85", X"7B", X"4C", X"AE", X"A7", X"8A", X"69", X"11", X"AA", X"9A", X"20", X"79", X"00", 
		X"C9", X"2C", X"D0", X"F1", X"20", X"73", X"00", X"20", X"24", X"AD", X"20", X"9E", X"AD", X"18", X"24", X"38", 
		X"24", X"0D", X"30", X"03", X"B0", X"03", X"60", X"B0", X"FD", X"A2", X"16", X"4C", X"37", X"A4", X"A6", X"7A", 
		X"D0", X"02", X"C6", X"7B", X"C6", X"7A", X"A2", X"00", X"24", X"48", X"8A", X"48", X"A9", X"01", X"20", X"FB", 
		X"A3", X"20", X"83", X"AE", X"A9", X"00", X"85", X"4D", X"20", X"79", X"00", X"38", X"E9", X"B1", X"90", X"17", 
		X"C9", X"03", X"B0", X"13", X"C9", X"01", X"2A", X"49", X"01", X"45", X"4D", X"C5", X"4D", X"90", X"61", X"85", 
		X"4D", X"20", X"73", X"00", X"4C", X"BB", X"AD", X"A6", X"4D", X"D0", X"2C", X"B0", X"7B", X"69", X"07", X"90", 
		X"77", X"65", X"0D", X"D0", X"03", X"4C", X"3D", X"B6", X"69", X"FF", X"85", X"22", X"0A", X"65", X"22", X"A8", 
		X"68", X"D9", X"80", X"A0", X"B0", X"67", X"20", X"8D", X"AD", X"48", X"20", X"20", X"AE", X"68", X"A4", X"4B", 
		X"10", X"17", X"AA", X"F0", X"56", X"D0", X"5F", X"46", X"0D", X"8A", X"2A", X"A6", X"7A", X"D0", X"02", X"C6", 
		X"7B", X"C6", X"7A", X"A0", X"1B", X"85", X"4D", X"D0", X"D7", X"D9", X"80", X"A0", X"B0", X"48", X"90", X"D9", 
		X"B9", X"82", X"A0", X"48", X"B9", X"81", X"A0", X"48", X"20", X"33", X"AE", X"A5", X"4D", X"4C", X"A9", X"AD", 
		X"4C", X"08", X"AF", X"A5", X"66", X"BE", X"80", X"A0", X"A8", X"68", X"85", X"22", X"E6", X"22", X"68", X"85", 
		X"23", X"98", X"48", X"20", X"1B", X"BC", X"A5", X"65", X"48", X"A5", X"64", X"48", X"A5", X"63", X"48", X"A5", 
		X"62", X"48", X"A5", X"61", X"48", X"6C", X"22", X"00", X"A0", X"FF", X"68", X"F0", X"23", X"C9", X"64", X"F0", 
		X"03", X"20", X"8D", X"AD", X"84", X"4B", X"68", X"4A", X"85", X"12", X"68", X"85", X"69", X"68", X"85", X"6A", 
		X"68", X"85", X"6B", X"68", X"85", X"6C", X"68", X"85", X"6D", X"68", X"85", X"6E", X"45", X"66", X"85", X"6F", 
		X"A5", X"61", X"60", X"6C", X"0A", X"03", X"A9", X"00", X"85", X"0D", X"20", X"73", X"00", X"B0", X"03", X"4C", 
		X"F3", X"BC", X"20", X"13", X"B1", X"90", X"03", X"4C", X"28", X"AF", X"C9", X"FF", X"D0", X"0F", X"A9", X"A8", 
		X"A0", X"AE", X"20", X"A2", X"BB", X"4C", X"73", X"00", X"82", X"49", X"0F", X"DA", X"A1", X"C9", X"2E", X"F0", 
		X"DE", X"C9", X"AB", X"F0", X"58", X"C9", X"AA", X"F0", X"D1", X"C9", X"22", X"D0", X"0F", X"A5", X"7A", X"A4", 
		X"7B", X"69", X"00", X"90", X"01", X"C8", X"20", X"87", X"B4", X"4C", X"E2", X"B7", X"C9", X"A8", X"D0", X"13", 
		X"A0", X"18", X"D0", X"3B", X"20", X"BF", X"B1", X"A5", X"65", X"49", X"FF", X"A8", X"A5", X"64", X"49", X"FF", 
		X"4C", X"91", X"B3", X"C9", X"A5", X"D0", X"03", X"4C", X"F4", X"B3", X"C9", X"B4", X"90", X"03", X"4C", X"A7", 
		X"AF", X"20", X"FA", X"AE", X"20", X"9E", X"AD", X"A9", X"29", X"2C", X"A9", X"28", X"2C", X"A9", X"2C", X"A0", 
		X"00", X"D1", X"7A", X"D0", X"03", X"4C", X"73", X"00", X"A2", X"0B", X"4C", X"37", X"A4", X"A0", X"15", X"68", 
		X"68", X"4C", X"FA", X"AD", X"38", X"A5", X"64", X"E9", X"00", X"A5", X"65", X"E9", X"A0", X"90", X"08", X"A9", 
		X"A2", X"E5", X"64", X"A9", X"E3", X"E5", X"65", X"60", X"20", X"8B", X"B0", X"85", X"64", X"84", X"65", X"A6", 
		X"45", X"A4", X"46", X"A5", X"0D", X"F0", X"26", X"A9", X"00", X"85", X"70", X"20", X"14", X"AF", X"90", X"1C", 
		X"E0", X"54", X"D0", X"18", X"C0", X"C9", X"D0", X"14", X"20", X"84", X"AF", X"84", X"5E", X"88", X"84", X"71", 
		X"A0", X"06", X"84", X"5D", X"A0", X"24", X"20", X"68", X"BE", X"4C", X"6F", X"B4", X"60", X"24", X"0E", X"10", 
		X"0D", X"A0", X"00", X"B1", X"64", X"AA", X"C8", X"B1", X"64", X"A8", X"8A", X"4C", X"91", X"B3", X"20", X"14", 
		X"AF", X"90", X"2D", X"E0", X"54", X"D0", X"1B", X"C0", X"49", X"D0", X"25", X"20", X"84", X"AF", X"98", X"A2", 
		X"A0", X"4C", X"4F", X"BC", X"20", X"DE", X"FF", X"86", X"64", X"84", X"63", X"85", X"65", X"A0", X"00", X"84", 
		X"62", X"60", X"E0", X"53", X"D0", X"0A", X"C0", X"54", X"D0", X"06", X"20", X"B7", X"FF", X"4C", X"3C", X"BC", 
		X"A5", X"64", X"A4", X"65", X"4C", X"A2", X"BB", X"0A", X"48", X"AA", X"20", X"73", X"00", X"E0", X"8F", X"90", 
		X"20", X"20", X"FA", X"AE", X"20", X"9E", X"AD", X"20", X"FD", X"AE", X"20", X"8F", X"AD", X"68", X"AA", X"A5", 
		X"65", X"48", X"A5", X"64", X"48", X"8A", X"48", X"20", X"9E", X"B7", X"68", X"A8", X"8A", X"48", X"4C", X"D6", 
		X"AF", X"20", X"F1", X"AE", X"68", X"A8", X"B9", X"EA", X"9F", X"85", X"55", X"B9", X"EB", X"9F", X"85", X"56", 
		X"20", X"54", X"00", X"4C", X"8D", X"AD", X"A0", X"FF", X"2C", X"A0", X"00", X"84", X"0B", X"20", X"BF", X"B1", 
		X"A5", X"64", X"45", X"0B", X"85", X"07", X"A5", X"65", X"45", X"0B", X"85", X"08", X"20", X"FC", X"BB", X"20", 
		X"BF", X"B1", X"A5", X"65", X"45", X"0B", X"25", X"08", X"45", X"0B", X"A8", X"A5", X"64", X"45", X"0B", X"25", 
		X"07", X"45", X"0B", X"4C", X"91", X"B3", X"20", X"90", X"AD", X"B0", X"13", X"A5", X"6E", X"09", X"7F", X"25", 
		X"6A", X"85", X"6A", X"A9", X"69", X"A0", X"00", X"20", X"5B", X"BC", X"AA", X"4C", X"61", X"B0", X"A9", X"00", 
		X"85", X"0D", X"C6", X"4D", X"20", X"A6", X"B6", X"85", X"61", X"86", X"62", X"84", X"63", X"A5", X"6C", X"A4", 
		X"6D", X"20", X"AA", X"B6", X"86", X"6C", X"84", X"6D", X"AA", X"38", X"E5", X"61", X"F0", X"08", X"A9", X"01", 
		X"90", X"04", X"A6", X"61", X"A9", X"FF", X"85", X"66", X"A0", X"FF", X"E8", X"C8", X"CA", X"D0", X"07", X"A6", 
		X"66", X"30", X"0F", X"18", X"90", X"0C", X"B1", X"6C", X"D1", X"62", X"F0", X"EF", X"A2", X"FF", X"B0", X"02", 
		X"A2", X"01", X"E8", X"8A", X"2A", X"25", X"12", X"F0", X"02", X"A9", X"FF", X"4C", X"3C", X"BC", X"20", X"FD", 
		X"AE", X"AA", X"20", X"90", X"B0", X"20", X"79", X"00", X"D0", X"F4", X"60", X"A2", X"00", X"20", X"79", X"00", 
		X"86", X"0C", X"85", X"45", X"20", X"79", X"00", X"20", X"13", X"B1", X"B0", X"03", X"4C", X"08", X"AF", X"A2", 
		X"00", X"86", X"0D", X"86", X"0E", X"20", X"73", X"00", X"90", X"05", X"20", X"13", X"B1", X"90", X"0B", X"AA", 
		X"20", X"73", X"00", X"90", X"FB", X"20", X"13", X"B1", X"B0", X"F6", X"C9", X"24", X"D0", X"06", X"A9", X"FF", 
		X"85", X"0D", X"D0", X"10", X"C9", X"25", X"D0", X"13", X"A5", X"10", X"D0", X"D0", X"A9", X"80", X"85", X"0E", 
		X"05", X"45", X"85", X"45", X"8A", X"09", X"80", X"AA", X"20", X"73", X"00", X"86", X"46", X"38", X"05", X"10", 
		X"E9", X"28", X"D0", X"03", X"4C", X"D1", X"B1", X"A0", X"00", X"84", X"10", X"A5", X"2D", X"A6", X"2E", X"86", 
		X"60", X"85", X"5F", X"E4", X"30", X"D0", X"04", X"C5", X"2F", X"F0", X"22", X"A5", X"45", X"D1", X"5F", X"D0", 
		X"08", X"A5", X"46", X"C8", X"D1", X"5F", X"F0", X"7D", X"88", X"18", X"A5", X"5F", X"69", X"07", X"90", X"E1", 
		X"E8", X"D0", X"DC", X"C9", X"41", X"90", X"05", X"E9", X"5B", X"38", X"E9", X"A5", X"60", X"68", X"48", X"C9", 
		X"2A", X"D0", X"05", X"A9", X"13", X"A0", X"BF", X"60", X"A5", X"45", X"A4", X"46", X"C9", X"54", X"D0", X"0B", 
		X"C0", X"C9", X"F0", X"EF", X"C0", X"49", X"D0", X"03", X"4C", X"08", X"AF", X"C9", X"53", X"D0", X"04", X"C0", 
		X"54", X"F0", X"F5", X"A5", X"2F", X"A4", X"30", X"85", X"5F", X"84", X"60", X"A5", X"31", X"A4", X"32", X"85", 
		X"5A", X"84", X"5B", X"18", X"69", X"07", X"90", X"01", X"C8", X"85", X"58", X"84", X"59", X"20", X"B8", X"A3", 
		X"A5", X"58", X"A4", X"59", X"C8", X"85", X"2F", X"84", X"30", X"A0", X"00", X"A5", X"45", X"91", X"5F", X"C8", 
		X"A5", X"46", X"91", X"5F", X"A9", X"00", X"C8", X"91", X"5F", X"C8", X"91", X"5F", X"C8", X"91", X"5F", X"C8", 
		X"91", X"5F", X"C8", X"91", X"5F", X"A5", X"5F", X"18", X"69", X"02", X"A4", X"60", X"90", X"01", X"C8", X"85", 
		X"47", X"84", X"48", X"60", X"A5", X"0B", X"0A", X"69", X"05", X"65", X"5F", X"A4", X"60", X"90", X"01", X"C8", 
		X"85", X"58", X"84", X"59", X"60", X"90", X"80", X"00", X"00", X"00", X"20", X"BF", X"B1", X"A5", X"64", X"A4", 
		X"65", X"60", X"20", X"73", X"00", X"20", X"9E", X"AD", X"20", X"8D", X"AD", X"A5", X"66", X"30", X"0D", X"A5", 
		X"61", X"C9", X"90", X"90", X"09", X"A9", X"A5", X"A0", X"B1", X"20", X"5B", X"BC", X"D0", X"7A", X"4C", X"9B", 
		X"BC", X"A5", X"0C", X"05", X"0E", X"48", X"A5", X"0D", X"48", X"A0", X"00", X"98", X"48", X"A5", X"46", X"48", 
		X"A5", X"45", X"48", X"20", X"B2", X"B1", X"68", X"85", X"45", X"68", X"85", X"46", X"68", X"A8", X"BA", X"BD", 
		X"02", X"01", X"48", X"BD", X"01", X"01", X"48", X"A5", X"64", X"9D", X"02", X"01", X"A5", X"65", X"9D", X"01", 
		X"01", X"C8", X"20", X"79", X"00", X"C9", X"2C", X"F0", X"D2", X"84", X"0B", X"20", X"F7", X"AE", X"68", X"85", 
		X"0D", X"68", X"85", X"0E", X"29", X"7F", X"85", X"0C", X"A6", X"2F", X"A5", X"30", X"86", X"5F", X"85", X"60", 
		X"C5", X"32", X"D0", X"04", X"E4", X"31", X"F0", X"39", X"A0", X"00", X"B1", X"5F", X"C8", X"C5", X"45", X"D0", 
		X"06", X"A5", X"46", X"D1", X"5F", X"F0", X"16", X"C8", X"B1", X"5F", X"18", X"65", X"5F", X"AA", X"C8", X"B1", 
		X"5F", X"65", X"60", X"90", X"D7", X"A2", X"12", X"2C", X"A2", X"0E", X"4C", X"37", X"A4", X"A2", X"13", X"A5", 
		X"0C", X"D0", X"F7", X"20", X"94", X"B1", X"A5", X"0B", X"A0", X"04", X"D1", X"5F", X"D0", X"E7", X"4C", X"EA", 
		X"B2", X"20", X"94", X"B1", X"20", X"08", X"A4", X"A0", X"00", X"84", X"72", X"A2", X"05", X"A5", X"45", X"91", 
		X"5F", X"10", X"01", X"CA", X"C8", X"A5", X"46", X"91", X"5F", X"10", X"02", X"CA", X"CA", X"86", X"71", X"A5", 
		X"0B", X"C8", X"C8", X"C8", X"91", X"5F", X"A2", X"0B", X"A9", X"00", X"24", X"0C", X"50", X"08", X"68", X"18", 
		X"69", X"01", X"AA", X"68", X"69", X"00", X"C8", X"91", X"5F", X"C8", X"8A", X"91", X"5F", X"20", X"4C", X"B3", 
		X"86", X"71", X"85", X"72", X"A4", X"22", X"C6", X"0B", X"D0", X"DC", X"65", X"59", X"B0", X"5D", X"85", X"59", 
		X"A8", X"8A", X"65", X"58", X"90", X"03", X"C8", X"F0", X"52", X"20", X"08", X"A4", X"85", X"31", X"84", X"32", 
		X"A9", X"00", X"E6", X"72", X"A4", X"71", X"F0", X"05", X"88", X"91", X"58", X"D0", X"FB", X"C6", X"59", X"C6", 
		X"72", X"D0", X"F5", X"E6", X"59", X"38", X"A5", X"31", X"E5", X"5F", X"A0", X"02", X"91", X"5F", X"A5", X"32", 
		X"C8", X"E5", X"60", X"91", X"5F", X"A5", X"0C", X"D0", X"62", X"C8", X"B1", X"5F", X"85", X"0B", X"A9", X"00", 
		X"85", X"71", X"85", X"72", X"C8", X"68", X"AA", X"85", X"64", X"68", X"85", X"65", X"D1", X"5F", X"90", X"0E", 
		X"D0", X"06", X"C8", X"8A", X"D1", X"5F", X"90", X"07", X"4C", X"45", X"B2", X"4C", X"35", X"A4", X"C8", X"A5", 
		X"72", X"05", X"71", X"18", X"F0", X"0A", X"20", X"4C", X"B3", X"8A", X"65", X"64", X"AA", X"98", X"A4", X"22", 
		X"65", X"65", X"86", X"71", X"C6", X"0B", X"D0", X"CA", X"85", X"72", X"A2", X"05", X"A5", X"45", X"10", X"01", 
		X"CA", X"A5", X"46", X"10", X"02", X"CA", X"CA", X"86", X"28", X"A9", X"00", X"20", X"55", X"B3", X"8A", X"65", 
		X"58", X"85", X"47", X"98", X"65", X"59", X"85", X"48", X"A8", X"A5", X"47", X"60", X"84", X"22", X"B1", X"5F", 
		X"85", X"28", X"88", X"B1", X"5F", X"85", X"29", X"A9", X"10", X"85", X"5D", X"A2", X"00", X"A0", X"00", X"8A", 
		X"0A", X"AA", X"98", X"2A", X"A8", X"B0", X"A4", X"06", X"71", X"26", X"72", X"90", X"0B", X"18", X"8A", X"65", 
		X"28", X"AA", X"98", X"65", X"29", X"A8", X"B0", X"93", X"C6", X"5D", X"D0", X"E3", X"60", X"A5", X"0D", X"F0", 
		X"03", X"20", X"A6", X"B6", X"20", X"26", X"B5", X"38", X"A5", X"33", X"E5", X"31", X"A8", X"A5", X"34", X"E5", 
		X"32", X"A2", X"00", X"86", X"0D", X"85", X"62", X"84", X"63", X"A2", X"90", X"4C", X"44", X"BC", X"38", X"20", 
		X"F0", X"FF", X"A9", X"00", X"F0", X"EB", X"A6", X"3A", X"E8", X"D0", X"A0", X"A2", X"15", X"2C", X"A2", X"1B", 
		X"4C", X"37", X"A4", X"20", X"E1", X"B3", X"20", X"A6", X"B3", X"20", X"FA", X"AE", X"A9", X"80", X"85", X"10", 
		X"20", X"8B", X"B0", X"20", X"8D", X"AD", X"20", X"F7", X"AE", X"A9", X"B2", X"20", X"FF", X"AE", X"48", X"A5", 
		X"48", X"48", X"A5", X"47", X"48", X"A5", X"7B", X"48", X"A5", X"7A", X"48", X"20", X"F8", X"A8", X"4C", X"4F", 
		X"B4", X"A9", X"A5", X"20", X"FF", X"AE", X"09", X"80", X"85", X"10", X"20", X"92", X"B0", X"85", X"4E", X"84", 
		X"4F", X"4C", X"8D", X"AD", X"20", X"E1", X"B3", X"A5", X"4F", X"48", X"A5", X"4E", X"48", X"20", X"F1", X"AE", 
		X"20", X"8D", X"AD", X"68", X"85", X"4E", X"68", X"85", X"4F", X"A0", X"02", X"B1", X"4E", X"85", X"47", X"AA", 
		X"C8", X"B1", X"4E", X"F0", X"99", X"85", X"48", X"C8", X"B1", X"47", X"48", X"88", X"10", X"FA", X"A4", X"48", 
		X"20", X"D4", X"BB", X"A5", X"7B", X"48", X"A5", X"7A", X"48", X"B1", X"4E", X"85", X"7A", X"C8", X"B1", X"4E", 
		X"85", X"7B", X"A5", X"48", X"48", X"A5", X"47", X"48", X"20", X"8A", X"AD", X"68", X"85", X"4E", X"68", X"85", 
		X"4F", X"20", X"79", X"00", X"F0", X"03", X"4C", X"08", X"AF", X"68", X"85", X"7A", X"68", X"85", X"7B", X"A0", 
		X"00", X"68", X"91", X"4E", X"68", X"C8", X"91", X"4E", X"68", X"C8", X"91", X"4E", X"68", X"C8", X"91", X"4E", 
		X"68", X"C8", X"91", X"4E", X"60", X"20", X"8D", X"AD", X"A0", X"00", X"20", X"DF", X"BD", X"68", X"68", X"A9", 
		X"FF", X"A0", X"00", X"F0", X"12", X"A6", X"64", X"A4", X"65", X"86", X"50", X"84", X"51", X"20", X"F4", X"B4", 
		X"86", X"62", X"84", X"63", X"85", X"61", X"60", X"A2", X"22", X"86", X"07", X"86", X"08", X"85", X"6F", X"84", 
		X"70", X"85", X"62", X"84", X"63", X"A0", X"FF", X"C8", X"B1", X"6F", X"F0", X"0C", X"C5", X"07", X"F0", X"04", 
		X"C5", X"08", X"D0", X"F3", X"C9", X"22", X"F0", X"01", X"18", X"84", X"61", X"98", X"65", X"6F", X"85", X"71", 
		X"A6", X"70", X"90", X"01", X"E8", X"86", X"72", X"A5", X"70", X"F0", X"04", X"C9", X"02", X"D0", X"0B", X"98", 
		X"20", X"75", X"B4", X"A6", X"6F", X"A4", X"70", X"20", X"88", X"B6", X"A6", X"16", X"E0", X"22", X"D0", X"05", 
		X"A2", X"19", X"4C", X"37", X"A4", X"A5", X"61", X"95", X"00", X"A5", X"62", X"95", X"01", X"A5", X"63", X"95", 
		X"02", X"A0", X"00", X"86", X"64", X"84", X"65", X"84", X"70", X"88", X"84", X"0D", X"86", X"17", X"E8", X"E8", 
		X"E8", X"86", X"16", X"60", X"46", X"0F", X"48", X"49", X"FF", X"38", X"65", X"33", X"A4", X"34", X"B0", X"01", 
		X"88", X"C4", X"32", X"90", X"11", X"D0", X"04", X"C5", X"31", X"90", X"0B", X"85", X"33", X"84", X"34", X"85", 
		X"35", X"84", X"36", X"AA", X"68", X"60", X"A2", X"10", X"A5", X"0F", X"30", X"B6", X"20", X"26", X"B5", X"A9", 
		X"80", X"85", X"0F", X"68", X"D0", X"D0", X"A6", X"37", X"A5", X"38", X"86", X"33", X"85", X"34", X"A0", X"00", 
		X"84", X"4F", X"84", X"4E", X"A5", X"31", X"A6", X"32", X"85", X"5F", X"86", X"60", X"A9", X"19", X"A2", X"00", 
		X"85", X"22", X"86", X"23", X"C5", X"16", X"F0", X"05", X"20", X"C7", X"B5", X"F0", X"F7", X"A9", X"07", X"85", 
		X"53", X"A5", X"2D", X"A6", X"2E", X"85", X"22", X"86", X"23", X"E4", X"30", X"D0", X"04", X"C5", X"2F", X"F0", 
		X"05", X"20", X"BD", X"B5", X"F0", X"F3", X"85", X"58", X"86", X"59", X"A9", X"03", X"85", X"53", X"A5", X"58", 
		X"A6", X"59", X"E4", X"32", X"D0", X"07", X"C5", X"31", X"D0", X"03", X"4C", X"06", X"B6", X"85", X"22", X"86", 
		X"23", X"A0", X"00", X"B1", X"22", X"AA", X"C8", X"B1", X"22", X"08", X"C8", X"B1", X"22", X"65", X"58", X"85", 
		X"58", X"C8", X"B1", X"22", X"65", X"59", X"85", X"59", X"28", X"10", X"D3", X"8A", X"30", X"D0", X"C8", X"B1", 
		X"22", X"A0", X"00", X"0A", X"69", X"05", X"65", X"22", X"85", X"22", X"90", X"02", X"E6", X"23", X"A6", X"23", 
		X"E4", X"59", X"D0", X"04", X"C5", X"58", X"F0", X"BA", X"20", X"C7", X"B5", X"F0", X"F3", X"B1", X"22", X"30", 
		X"35", X"C8", X"B1", X"22", X"10", X"30", X"C8", X"B1", X"22", X"F0", X"2B", X"C8", X"B1", X"22", X"AA", X"C8", 
		X"B1", X"22", X"C5", X"34", X"90", X"06", X"D0", X"1E", X"E4", X"33", X"B0", X"1A", X"C5", X"60", X"90", X"16", 
		X"D0", X"04", X"E4", X"5F", X"90", X"10", X"86", X"5F", X"85", X"60", X"A5", X"22", X"A6", X"23", X"85", X"4E", 
		X"86", X"4F", X"A5", X"53", X"85", X"55", X"A5", X"53", X"18", X"65", X"22", X"85", X"22", X"90", X"02", X"E6", 
		X"23", X"A6", X"23", X"A0", X"00", X"60", X"A5", X"4F", X"05", X"4E", X"F0", X"F5", X"A5", X"55", X"29", X"04", 
		X"4A", X"A8", X"85", X"55", X"B1", X"4E", X"65", X"5F", X"85", X"5A", X"A5", X"60", X"69", X"00", X"85", X"5B", 
		X"A5", X"33", X"A6", X"34", X"85", X"58", X"86", X"59", X"20", X"BF", X"A3", X"A4", X"55", X"C8", X"A5", X"58", 
		X"91", X"4E", X"AA", X"E6", X"59", X"A5", X"59", X"C8", X"91", X"4E", X"4C", X"2A", X"B5", X"A5", X"65", X"48", 
		X"A5", X"64", X"48", X"20", X"83", X"AE", X"20", X"8F", X"AD", X"68", X"85", X"6F", X"68", X"85", X"70", X"A0", 
		X"00", X"B1", X"6F", X"18", X"71", X"64", X"90", X"05", X"A2", X"17", X"4C", X"37", X"A4", X"20", X"75", X"B4", 
		X"20", X"7A", X"B6", X"A5", X"50", X"A4", X"51", X"20", X"AA", X"B6", X"20", X"8C", X"B6", X"A5", X"6F", X"A4", 
		X"70", X"20", X"AA", X"B6", X"20", X"CA", X"B4", X"4C", X"B8", X"AD", X"A0", X"00", X"B1", X"6F", X"48", X"C8", 
		X"B1", X"6F", X"AA", X"C8", X"B1", X"6F", X"A8", X"68", X"86", X"22", X"84", X"23", X"A8", X"F0", X"0A", X"48", 
		X"88", X"B1", X"22", X"91", X"35", X"98", X"D0", X"F8", X"68", X"18", X"65", X"35", X"85", X"35", X"90", X"02", 
		X"E6", X"36", X"60", X"20", X"8F", X"AD", X"A5", X"64", X"A4", X"65", X"85", X"22", X"84", X"23", X"20", X"DB", 
		X"B6", X"08", X"A0", X"00", X"B1", X"22", X"48", X"C8", X"B1", X"22", X"AA", X"C8", X"B1", X"22", X"A8", X"68", 
		X"28", X"D0", X"13", X"C4", X"34", X"D0", X"0F", X"E4", X"33", X"D0", X"0B", X"48", X"18", X"65", X"33", X"85", 
		X"33", X"90", X"02", X"E6", X"34", X"68", X"86", X"22", X"84", X"23", X"60", X"C4", X"18", X"D0", X"0C", X"C5", 
		X"17", X"D0", X"08", X"85", X"16", X"E9", X"03", X"85", X"17", X"A0", X"00", X"60", X"20", X"A1", X"B7", X"8A", 
		X"48", X"A9", X"01", X"20", X"7D", X"B4", X"68", X"A0", X"00", X"91", X"62", X"68", X"68", X"4C", X"CA", X"B4", 
		X"20", X"61", X"B7", X"D1", X"50", X"98", X"90", X"04", X"B1", X"50", X"AA", X"98", X"48", X"8A", X"48", X"20", 
		X"7D", X"B4", X"A5", X"50", X"A4", X"51", X"20", X"AA", X"B6", X"68", X"A8", X"68", X"18", X"65", X"22", X"85", 
		X"22", X"90", X"02", X"E6", X"23", X"98", X"20", X"8C", X"B6", X"4C", X"CA", X"B4", X"20", X"61", X"B7", X"18", 
		X"F1", X"50", X"49", X"FF", X"4C", X"06", X"B7", X"A9", X"FF", X"85", X"65", X"20", X"79", X"00", X"C9", X"29", 
		X"F0", X"06", X"20", X"FD", X"AE", X"20", X"9E", X"B7", X"20", X"61", X"B7", X"F0", X"4B", X"CA", X"8A", X"48", 
		X"18", X"A2", X"00", X"F1", X"50", X"B0", X"B6", X"49", X"FF", X"C5", X"65", X"90", X"B1", X"A5", X"65", X"B0", 
		X"AD", X"20", X"F7", X"AE", X"68", X"A8", X"68", X"85", X"55", X"68", X"68", X"68", X"AA", X"68", X"85", X"50", 
		X"68", X"85", X"51", X"A5", X"55", X"48", X"98", X"48", X"A0", X"00", X"8A", X"60", X"20", X"82", X"B7", X"4C", 
		X"A2", X"B3", X"20", X"A3", X"B6", X"A2", X"00", X"86", X"0D", X"A8", X"60", X"20", X"82", X"B7", X"F0", X"08", 
		X"A0", X"00", X"B1", X"22", X"A8", X"4C", X"A2", X"B3", X"4C", X"48", X"B2", X"20", X"73", X"00", X"20", X"8A", 
		X"AD", X"20", X"B8", X"B1", X"A6", X"64", X"D0", X"F0", X"A6", X"65", X"4C", X"79", X"00", X"20", X"82", X"B7", 
		X"D0", X"03", X"4C", X"F7", X"B8", X"A6", X"7A", X"A4", X"7B", X"86", X"71", X"84", X"72", X"A6", X"22", X"86", 
		X"7A", X"18", X"65", X"22", X"85", X"24", X"A6", X"23", X"86", X"7B", X"90", X"01", X"E8", X"86", X"25", X"A0", 
		X"00", X"B1", X"24", X"48", X"98", X"91", X"24", X"20", X"79", X"00", X"20", X"F3", X"BC", X"68", X"A0", X"00", 
		X"91", X"24", X"A6", X"71", X"A4", X"72", X"86", X"7A", X"84", X"7B", X"60", X"20", X"8A", X"AD", X"20", X"F7", 
		X"B7", X"20", X"FD", X"AE", X"4C", X"9E", X"B7", X"A5", X"66", X"30", X"9D", X"A5", X"61", X"C9", X"91", X"B0", 
		X"97", X"20", X"9B", X"BC", X"A5", X"64", X"A4", X"65", X"84", X"14", X"85", X"15", X"60", X"A5", X"15", X"48", 
		X"A5", X"14", X"48", X"20", X"F7", X"B7", X"A0", X"00", X"B1", X"14", X"A8", X"68", X"85", X"14", X"68", X"85", 
		X"15", X"4C", X"A2", X"B3", X"20", X"EB", X"B7", X"8A", X"A0", X"00", X"91", X"14", X"60", X"20", X"EB", X"B7", 
		X"86", X"49", X"A2", X"00", X"20", X"79", X"00", X"F0", X"03", X"20", X"F1", X"B7", X"86", X"4A", X"A0", X"00", 
		X"B1", X"14", X"45", X"4A", X"25", X"49", X"F0", X"F8", X"60", X"A9", X"11", X"A0", X"BF", X"4C", X"67", X"B8", 
		X"20", X"8C", X"BA", X"A5", X"66", X"49", X"FF", X"85", X"66", X"45", X"6E", X"85", X"6F", X"A5", X"61", X"4C", 
		X"6A", X"B8", X"20", X"99", X"B9", X"90", X"3C", X"20", X"8C", X"BA", X"D0", X"03", X"4C", X"FC", X"BB", X"A6", 
		X"70", X"86", X"56", X"A2", X"69", X"A5", X"69", X"A8", X"F0", X"CE", X"38", X"E5", X"61", X"F0", X"24", X"90", 
		X"12", X"84", X"61", X"A4", X"6E", X"84", X"66", X"49", X"FF", X"69", X"00", X"A0", X"00", X"84", X"56", X"A2", 
		X"61", X"D0", X"04", X"A0", X"00", X"84", X"70", X"C9", X"F9", X"30", X"C7", X"A8", X"A5", X"70", X"56", X"01", 
		X"20", X"B0", X"B9", X"24", X"6F", X"10", X"57", X"A0", X"61", X"E0", X"69", X"F0", X"02", X"A0", X"69", X"38", 
		X"49", X"FF", X"65", X"56", X"85", X"70", X"B9", X"04", X"00", X"F5", X"04", X"85", X"65", X"B9", X"03", X"00", 
		X"F5", X"03", X"85", X"64", X"B9", X"02", X"00", X"F5", X"02", X"85", X"63", X"B9", X"01", X"00", X"F5", X"01", 
		X"85", X"62", X"B0", X"03", X"20", X"47", X"B9", X"A0", X"00", X"98", X"18", X"A6", X"62", X"D0", X"4A", X"A6", 
		X"63", X"86", X"62", X"A6", X"64", X"86", X"63", X"A6", X"65", X"86", X"64", X"A6", X"70", X"86", X"65", X"84", 
		X"70", X"69", X"08", X"C9", X"20", X"D0", X"E4", X"A9", X"00", X"85", X"61", X"85", X"66", X"60", X"65", X"56", 
		X"85", X"70", X"A5", X"65", X"65", X"6D", X"85", X"65", X"A5", X"64", X"65", X"6C", X"85", X"64", X"A5", X"63", 
		X"65", X"6B", X"85", X"63", X"A5", X"62", X"65", X"6A", X"85", X"62", X"4C", X"36", X"B9", X"69", X"01", X"06", 
		X"70", X"26", X"65", X"26", X"64", X"26", X"63", X"26", X"62", X"10", X"F2", X"38", X"E5", X"61", X"B0", X"C7", 
		X"49", X"FF", X"69", X"01", X"85", X"61", X"90", X"0E", X"E6", X"61", X"F0", X"42", X"66", X"62", X"66", X"63", 
		X"66", X"64", X"66", X"65", X"66", X"70", X"60", X"A5", X"66", X"49", X"FF", X"85", X"66", X"A5", X"62", X"49", 
		X"FF", X"85", X"62", X"A5", X"63", X"49", X"FF", X"85", X"63", X"A5", X"64", X"49", X"FF", X"85", X"64", X"A5", 
		X"65", X"49", X"FF", X"85", X"65", X"A5", X"70", X"49", X"FF", X"85", X"70", X"E6", X"70", X"D0", X"0E", X"E6", 
		X"65", X"D0", X"0A", X"E6", X"64", X"D0", X"06", X"E6", X"63", X"D0", X"02", X"E6", X"62", X"60", X"A2", X"0F", 
		X"4C", X"37", X"A4", X"A2", X"25", X"B4", X"04", X"84", X"70", X"B4", X"03", X"94", X"04", X"B4", X"02", X"94", 
		X"03", X"B4", X"01", X"94", X"02", X"A4", X"68", X"94", X"01", X"69", X"08", X"30", X"E8", X"F0", X"E6", X"E9", 
		X"08", X"A8", X"A5", X"70", X"B0", X"14", X"16", X"01", X"90", X"02", X"F6", X"01", X"76", X"01", X"76", X"01", 
		X"76", X"02", X"76", X"03", X"76", X"04", X"6A", X"C8", X"D0", X"EC", X"18", X"60", X"81", X"00", X"00", X"00", 
		X"00", X"03", X"7F", X"5E", X"56", X"CB", X"79", X"80", X"13", X"9B", X"0B", X"64", X"80", X"76", X"38", X"93", 
		X"16", X"82", X"38", X"AA", X"3B", X"20", X"80", X"35", X"04", X"F3", X"34", X"81", X"35", X"04", X"F3", X"34", 
		X"80", X"80", X"00", X"00", X"00", X"80", X"31", X"72", X"17", X"F8", X"20", X"2B", X"BC", X"F0", X"02", X"10", 
		X"03", X"4C", X"48", X"B2", X"A5", X"61", X"E9", X"7F", X"48", X"A9", X"80", X"85", X"61", X"A9", X"D6", X"A0", 
		X"B9", X"20", X"67", X"B8", X"A9", X"DB", X"A0", X"B9", X"20", X"0F", X"BB", X"A9", X"BC", X"A0", X"B9", X"20", 
		X"50", X"B8", X"A9", X"C1", X"A0", X"B9", X"20", X"43", X"E0", X"A9", X"E0", X"A0", X"B9", X"20", X"67", X"B8", 
		X"68", X"20", X"7E", X"BD", X"A9", X"E5", X"A0", X"B9", X"20", X"8C", X"BA", X"D0", X"03", X"4C", X"8B", X"BA", 
		X"20", X"B7", X"BA", X"A9", X"00", X"85", X"26", X"85", X"27", X"85", X"28", X"85", X"29", X"A5", X"70", X"20", 
		X"59", X"BA", X"A5", X"65", X"20", X"59", X"BA", X"A5", X"64", X"20", X"59", X"BA", X"A5", X"63", X"20", X"59", 
		X"BA", X"A5", X"62", X"20", X"5E", X"BA", X"4C", X"8F", X"BB", X"D0", X"03", X"4C", X"83", X"B9", X"4A", X"09", 
		X"80", X"A8", X"90", X"19", X"18", X"A5", X"29", X"65", X"6D", X"85", X"29", X"A5", X"28", X"65", X"6C", X"85", 
		X"28", X"A5", X"27", X"65", X"6B", X"85", X"27", X"A5", X"26", X"65", X"6A", X"85", X"26", X"66", X"26", X"66", 
		X"27", X"66", X"28", X"66", X"29", X"66", X"70", X"98", X"4A", X"D0", X"D6", X"60", X"85", X"22", X"84", X"23", 
		X"A0", X"04", X"B1", X"22", X"85", X"6D", X"88", X"B1", X"22", X"85", X"6C", X"88", X"B1", X"22", X"85", X"6B", 
		X"88", X"B1", X"22", X"85", X"6E", X"45", X"66", X"85", X"6F", X"A5", X"6E", X"09", X"80", X"85", X"6A", X"88", 
		X"B1", X"22", X"85", X"69", X"A5", X"61", X"60", X"A5", X"69", X"F0", X"1F", X"18", X"65", X"61", X"90", X"04", 
		X"30", X"1D", X"18", X"2C", X"10", X"14", X"69", X"80", X"85", X"61", X"D0", X"03", X"4C", X"FB", X"B8", X"A5", 
		X"6F", X"85", X"66", X"60", X"A5", X"66", X"49", X"FF", X"30", X"05", X"68", X"68", X"4C", X"F7", X"B8", X"4C", 
		X"7E", X"B9", X"20", X"0C", X"BC", X"AA", X"F0", X"10", X"18", X"69", X"02", X"B0", X"F2", X"A2", X"00", X"86", 
		X"6F", X"20", X"77", X"B8", X"E6", X"61", X"F0", X"E7", X"60", X"84", X"20", X"00", X"00", X"00", X"20", X"0C", 
		X"BC", X"A9", X"F9", X"A0", X"BA", X"A2", X"00", X"86", X"6F", X"20", X"A2", X"BB", X"4C", X"12", X"BB", X"20", 
		X"8C", X"BA", X"F0", X"76", X"20", X"1B", X"BC", X"A9", X"00", X"38", X"E5", X"61", X"85", X"61", X"20", X"B7", 
		X"BA", X"E6", X"61", X"F0", X"BA", X"A2", X"FC", X"A9", X"01", X"A4", X"6A", X"C4", X"62", X"D0", X"10", X"A4", 
		X"6B", X"C4", X"63", X"D0", X"0A", X"A4", X"6C", X"C4", X"64", X"D0", X"04", X"A4", X"6D", X"C4", X"65", X"08", 
		X"2A", X"90", X"09", X"E8", X"95", X"29", X"F0", X"32", X"10", X"34", X"A9", X"01", X"28", X"B0", X"0E", X"06", 
		X"6D", X"26", X"6C", X"26", X"6B", X"26", X"6A", X"B0", X"E6", X"30", X"CE", X"10", X"E2", X"A8", X"A5", X"6D", 
		X"E5", X"65", X"85", X"6D", X"A5", X"6C", X"E5", X"64", X"85", X"6C", X"A5", X"6B", X"E5", X"63", X"85", X"6B", 
		X"A5", X"6A", X"E5", X"62", X"85", X"6A", X"98", X"4C", X"4F", X"BB", X"A9", X"40", X"D0", X"CE", X"0A", X"0A", 
		X"0A", X"0A", X"0A", X"0A", X"85", X"70", X"28", X"4C", X"8F", X"BB", X"A2", X"14", X"4C", X"37", X"A4", X"A5", 
		X"26", X"85", X"62", X"A5", X"27", X"85", X"63", X"A5", X"28", X"85", X"64", X"A5", X"29", X"85", X"65", X"4C", 
		X"D7", X"B8", X"85", X"22", X"84", X"23", X"A0", X"04", X"B1", X"22", X"85", X"65", X"88", X"B1", X"22", X"85", 
		X"64", X"88", X"B1", X"22", X"85", X"63", X"88", X"B1", X"22", X"85", X"66", X"09", X"80", X"85", X"62", X"88", 
		X"B1", X"22", X"85", X"61", X"84", X"70", X"60", X"A2", X"5C", X"2C", X"A2", X"57", X"A0", X"00", X"F0", X"04", 
		X"A6", X"49", X"A4", X"4A", X"20", X"1B", X"BC", X"86", X"22", X"84", X"23", X"A0", X"04", X"A5", X"65", X"91", 
		X"22", X"88", X"A5", X"64", X"91", X"22", X"88", X"A5", X"63", X"91", X"22", X"88", X"A5", X"66", X"09", X"7F", 
		X"25", X"62", X"91", X"22", X"88", X"A5", X"61", X"91", X"22", X"84", X"70", X"60", X"A5", X"6E", X"85", X"66", 
		X"A2", X"05", X"B5", X"68", X"95", X"60", X"CA", X"D0", X"F9", X"86", X"70", X"60", X"20", X"1B", X"BC", X"A2", 
		X"06", X"B5", X"60", X"95", X"68", X"CA", X"D0", X"F9", X"86", X"70", X"60", X"A5", X"61", X"F0", X"FB", X"06", 
		X"70", X"90", X"F7", X"20", X"6F", X"B9", X"D0", X"F2", X"4C", X"38", X"B9", X"A5", X"61", X"F0", X"09", X"A5", 
		X"66", X"2A", X"A9", X"FF", X"B0", X"02", X"A9", X"01", X"60", X"20", X"2B", X"BC", X"85", X"62", X"A9", X"00", 
		X"85", X"63", X"A2", X"88", X"A5", X"62", X"49", X"FF", X"2A", X"A9", X"00", X"85", X"65", X"85", X"64", X"86", 
		X"61", X"85", X"70", X"85", X"66", X"4C", X"D2", X"B8", X"46", X"66", X"60", X"85", X"24", X"84", X"25", X"A0", 
		X"00", X"B1", X"24", X"C8", X"AA", X"F0", X"C4", X"B1", X"24", X"45", X"66", X"30", X"C2", X"E4", X"61", X"D0", 
		X"21", X"B1", X"24", X"09", X"80", X"C5", X"62", X"D0", X"19", X"C8", X"B1", X"24", X"C5", X"63", X"D0", X"12", 
		X"C8", X"B1", X"24", X"C5", X"64", X"D0", X"0B", X"C8", X"A9", X"7F", X"C5", X"70", X"B1", X"24", X"E5", X"65", 
		X"F0", X"28", X"A5", X"66", X"90", X"02", X"49", X"FF", X"4C", X"31", X"BC", X"A5", X"61", X"F0", X"4A", X"38", 
		X"E9", X"A0", X"24", X"66", X"10", X"09", X"AA", X"A9", X"FF", X"85", X"68", X"20", X"4D", X"B9", X"8A", X"A2", 
		X"61", X"C9", X"F9", X"10", X"06", X"20", X"99", X"B9", X"84", X"68", X"60", X"A8", X"A5", X"66", X"29", X"80", 
		X"46", X"62", X"05", X"62", X"85", X"62", X"20", X"B0", X"B9", X"84", X"68", X"60", X"A5", X"61", X"C9", X"A0", 
		X"B0", X"20", X"20", X"9B", X"BC", X"84", X"70", X"A5", X"66", X"84", X"66", X"49", X"80", X"2A", X"A9", X"A0", 
		X"85", X"61", X"A5", X"65", X"85", X"07", X"4C", X"D2", X"B8", X"85", X"62", X"85", X"63", X"85", X"64", X"85", 
		X"65", X"A8", X"60", X"A0", X"00", X"A2", X"0A", X"94", X"5D", X"CA", X"10", X"FB", X"90", X"0F", X"C9", X"2D", 
		X"D0", X"04", X"86", X"67", X"F0", X"04", X"C9", X"2B", X"D0", X"05", X"20", X"73", X"00", X"90", X"5B", X"C9", 
		X"2E", X"F0", X"2E", X"C9", X"45", X"D0", X"30", X"20", X"73", X"00", X"90", X"17", X"C9", X"AB", X"F0", X"0E", 
		X"C9", X"2D", X"F0", X"0A", X"C9", X"AA", X"F0", X"08", X"C9", X"2B", X"F0", X"04", X"D0", X"07", X"66", X"60", 
		X"20", X"73", X"00", X"90", X"5C", X"24", X"60", X"10", X"0E", X"A9", X"00", X"38", X"E5", X"5E", X"4C", X"49", 
		X"BD", X"66", X"5F", X"24", X"5F", X"50", X"C3", X"A5", X"5E", X"38", X"E5", X"5D", X"85", X"5E", X"F0", X"12", 
		X"10", X"09", X"20", X"FE", X"BA", X"E6", X"5E", X"D0", X"F9", X"F0", X"07", X"20", X"E2", X"BA", X"C6", X"5E", 
		X"D0", X"F9", X"A5", X"67", X"30", X"01", X"60", X"4C", X"B4", X"BF", X"48", X"24", X"5F", X"10", X"02", X"E6", 
		X"5D", X"20", X"E2", X"BA", X"68", X"38", X"E9", X"30", X"20", X"7E", X"BD", X"4C", X"0A", X"BD", X"48", X"20", 
		X"0C", X"BC", X"68", X"20", X"3C", X"BC", X"A5", X"6E", X"45", X"66", X"85", X"6F", X"A6", X"61", X"4C", X"6A", 
		X"B8", X"A5", X"5E", X"C9", X"0A", X"90", X"09", X"A9", X"64", X"24", X"60", X"30", X"11", X"4C", X"7E", X"B9", 
		X"0A", X"0A", X"18", X"65", X"5E", X"0A", X"18", X"A0", X"00", X"71", X"7A", X"38", X"E9", X"30", X"85", X"5E", 
		X"4C", X"30", X"BD", X"9B", X"3E", X"BC", X"1F", X"FD", X"9E", X"6E", X"6B", X"27", X"FD", X"9E", X"6E", X"6B", 
		X"28", X"00", X"A9", X"71", X"A0", X"A3", X"20", X"DA", X"BD", X"A5", X"3A", X"A6", X"39", X"85", X"62", X"86", 
		X"63", X"A2", X"90", X"38", X"20", X"49", X"BC", X"20", X"DF", X"BD", X"4C", X"1E", X"AB", X"A0", X"01", X"A9", 
		X"20", X"24", X"66", X"10", X"02", X"A9", X"2D", X"99", X"FF", X"00", X"85", X"66", X"84", X"71", X"C8", X"A9", 
		X"30", X"A6", X"61", X"D0", X"03", X"4C", X"04", X"BF", X"A9", X"00", X"E0", X"80", X"F0", X"02", X"B0", X"09", 
		X"A9", X"BD", X"A0", X"BD", X"20", X"28", X"BA", X"A9", X"F7", X"85", X"5D", X"A9", X"B8", X"A0", X"BD", X"20", 
		X"5B", X"BC", X"F0", X"1E", X"10", X"12", X"A9", X"B3", X"A0", X"BD", X"20", X"5B", X"BC", X"F0", X"02", X"10", 
		X"0E", X"20", X"E2", X"BA", X"C6", X"5D", X"D0", X"EE", X"20", X"FE", X"BA", X"E6", X"5D", X"D0", X"DC", X"20", 
		X"49", X"B8", X"20", X"9B", X"BC", X"A2", X"01", X"A5", X"5D", X"18", X"69", X"0A", X"30", X"09", X"C9", X"0B", 
		X"B0", X"06", X"69", X"FF", X"AA", X"A9", X"02", X"38", X"E9", X"02", X"85", X"5E", X"86", X"5D", X"8A", X"F0", 
		X"02", X"10", X"13", X"A4", X"71", X"A9", X"2E", X"C8", X"99", X"FF", X"00", X"8A", X"F0", X"06", X"A9", X"30", 
		X"C8", X"99", X"FF", X"00", X"84", X"71", X"A0", X"00", X"A2", X"80", X"A5", X"65", X"18", X"79", X"19", X"BF", 
		X"85", X"65", X"A5", X"64", X"79", X"18", X"BF", X"85", X"64", X"A5", X"63", X"79", X"17", X"BF", X"85", X"63", 
		X"A5", X"62", X"79", X"16", X"BF", X"85", X"62", X"E8", X"B0", X"04", X"10", X"DE", X"30", X"02", X"30", X"DA", 
		X"8A", X"90", X"04", X"49", X"FF", X"69", X"0A", X"69", X"2F", X"C8", X"C8", X"C8", X"C8", X"84", X"47", X"A4", 
		X"71", X"C8", X"AA", X"29", X"7F", X"99", X"FF", X"00", X"C6", X"5D", X"D0", X"06", X"A9", X"2E", X"C8", X"99", 
		X"FF", X"00", X"84", X"71", X"A4", X"47", X"8A", X"49", X"FF", X"29", X"80", X"AA", X"C0", X"24", X"F0", X"04", 
		X"C0", X"3C", X"D0", X"A6", X"A4", X"71", X"B9", X"FF", X"00", X"88", X"C9", X"30", X"F0", X"F8", X"C9", X"2E", 
		X"F0", X"01", X"C8", X"A9", X"2B", X"A6", X"5E", X"F0", X"2E", X"10", X"08", X"A9", X"00", X"38", X"E5", X"5E", 
		X"AA", X"A9", X"2D", X"99", X"01", X"01", X"A9", X"45", X"99", X"00", X"01", X"8A", X"A2", X"2F", X"38", X"E8", 
		X"E9", X"0A", X"B0", X"FB", X"69", X"3A", X"99", X"03", X"01", X"8A", X"99", X"02", X"01", X"A9", X"00", X"99", 
		X"04", X"01", X"F0", X"08", X"99", X"FF", X"00", X"A9", X"00", X"99", X"00", X"01", X"A9", X"00", X"A0", X"01", 
		X"60", X"80", X"00", X"00", X"00", X"00", X"FA", X"0A", X"1F", X"00", X"00", X"98", X"96", X"80", X"FF", X"F0", 
		X"BD", X"C0", X"00", X"01", X"86", X"A0", X"FF", X"FF", X"D8", X"F0", X"00", X"00", X"03", X"E8", X"FF", X"FF", 
		X"FF", X"9C", X"00", X"00", X"00", X"0A", X"FF", X"FF", X"FF", X"FF", X"FF", X"DF", X"0A", X"80", X"00", X"03", 
		X"4B", X"C0", X"FF", X"FF", X"73", X"60", X"00", X"00", X"0E", X"10", X"FF", X"FF", X"FD", X"A8", X"00", X"00", 
		X"00", X"3C", X"EC", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", 
		X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", 
		X"AA", X"20", X"0C", X"BC", X"A9", X"11", X"A0", X"BF", X"20", X"A2", X"BB", X"F0", X"70", X"A5", X"69", X"D0", 
		X"03", X"4C", X"F9", X"B8", X"A2", X"4E", X"A0", X"00", X"20", X"D4", X"BB", X"A5", X"6E", X"10", X"0F", X"20", 
		X"CC", X"BC", X"A9", X"4E", X"A0", X"00", X"20", X"5B", X"BC", X"D0", X"03", X"98", X"A4", X"07", X"20", X"FE", 
		X"BB", X"98", X"48", X"20", X"EA", X"B9", X"A9", X"4E", X"A0", X"00", X"20", X"28", X"BA", X"20", X"ED", X"BF", 
		X"68", X"4A", X"90", X"0A", X"A5", X"61", X"F0", X"06", X"A5", X"66", X"49", X"FF", X"85", X"66", X"60", X"81", 
		X"38", X"AA", X"3B", X"29", X"07", X"71", X"34", X"58", X"3E", X"56", X"74", X"16", X"7E", X"B3", X"1B", X"77", 
		X"2F", X"EE", X"E3", X"85", X"7A", X"1D", X"84", X"1C", X"2A", X"7C", X"63", X"59", X"58", X"0A", X"7E", X"75", 
		X"FD", X"E7", X"C6", X"80", X"31", X"72", X"18", X"10", X"81", X"00", X"00", X"00", X"00", X"A9", X"BF", X"A0", 
		X"BF", X"20", X"28", X"BA", X"A5", X"70", X"69", X"50", X"90", X"03", X"20", X"23", X"BC", X"4C", X"00", X"E0" 
	);
--	signal localAddr : unsigned(11 downto 0);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			do <= romData(to_integer(addr)) after 2 ns;
		end if;
	end process;
end Behavioral;

